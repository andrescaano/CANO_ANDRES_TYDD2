library verilog;
use verilog.vl_types.all;
entity Parte_B_vlg_vec_tst is
end Parte_B_vlg_vec_tst;

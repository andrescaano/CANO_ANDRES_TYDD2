library verilog;
use verilog.vl_types.all;
entity Parte_D_vlg_check_tst is
    port(
        z               : in     vl_logic_vector(0 to 3);
        sampler_rx      : in     vl_logic
    );
end Parte_D_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Ej1_Cano_vlg_vec_tst is
end Ej1_Cano_vlg_vec_tst;

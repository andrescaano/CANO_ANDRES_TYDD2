library verilog;
use verilog.vl_types.all;
entity Template_vlg_vec_tst is
end Template_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Ej1_Cano_vlg_check_tst is
    port(
        LED             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Ej1_Cano_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Ej1_Cano is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        LED             : out    vl_logic
    );
end Ej1_Cano;

library verilog;
use verilog.vl_types.all;
entity Parte_B_vlg_check_tst is
    port(
        output_Cout     : in     vl_logic;
        output_S        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Parte_B_vlg_check_tst;
